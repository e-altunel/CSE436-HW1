* SPICE3 file created from /output/not/not.ext - technology: scmos

.option scale=0.12u

M1000 y a gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1001 y a vdd vdd pfet w=8 l=2
+  ad=40 pd=26 as=40 ps=26
