* SPICE3 file created from /output/nor/nor.ext - technology: scmos

.option scale=0.12u

M1000 gnd a y Gnd nfet w=4 l=2
+  ad=24 pd=20 as=40 ps=36
M1001 y b a_11_81# vdd pfet w=8 l=2
+  ad=40 pd=26 as=48 ps=28
M1002 y b gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_11_81# a vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
